* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlclkp_2 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_27_74# a_83_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VPWR a_1041_387# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_1044_119# a_27_74# a_1041_387# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_315_48# a_315_338# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X4 a_508_508# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X5 a_494_118# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_1041_387# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 VGND a_1041_387# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 GCLK a_1041_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 a_83_244# a_315_338# a_494_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 VGND CLK a_1044_119# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_315_48# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR GATE a_264_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X13 a_83_244# a_315_48# a_508_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 a_267_74# a_315_48# a_83_244# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 VGND a_315_48# a_315_338# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_315_48# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X17 GCLK a_1041_387# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VGND GATE a_267_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_27_74# a_83_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_264_392# a_315_338# a_83_244# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X21 VPWR CLK a_1041_387# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
