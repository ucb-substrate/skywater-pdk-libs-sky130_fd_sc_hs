* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_851_368# A3 a_762_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VPWR a_110_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VPWR B1 a_110_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X3 a_1213_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 VPWR a_110_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 VGND A3 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_851_368# A4 a_110_48# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VGND a_110_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_523_124# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_523_124# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 VGND A2 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VGND A1 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_762_368# A2 a_1213_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_523_124# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 X a_110_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 X a_110_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 X a_110_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_110_48# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X18 X a_110_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 VPWR A1 a_1213_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 a_762_368# A3 a_851_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_523_124# B1 a_110_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 a_110_48# B1 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 VGND A4 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 a_523_124# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X25 a_1213_368# A2 a_762_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 a_110_48# A4 a_851_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 VGND a_110_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
