* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nand3b_2 A_N B C VGND VNB VPB VPWR Y
X0 Y a_27_94# a_403_54# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_403_54# B a_206_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_27_94# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 a_206_74# B a_403_54# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND C a_206_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 a_27_94# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_206_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_403_54# a_27_94# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 Y a_27_94# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_27_94# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
