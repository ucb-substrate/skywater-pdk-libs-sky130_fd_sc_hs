* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__xor3_1 A B C VGND VNB VPB VPWR X
X0 a_27_134# B a_384_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_452_288# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_416_86# a_452_288# a_27_134# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_27_134# B a_416_86# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X4 a_452_288# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_1215_396# C a_384_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 a_84_108# B a_416_86# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 VGND a_1215_396# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND A a_84_108# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_84_108# B a_384_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 a_416_86# a_1157_298# a_1215_396# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X11 a_384_392# a_452_288# a_27_134# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X12 a_384_392# a_1157_298# a_1215_396# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 VPWR a_1215_396# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_384_392# a_452_288# a_84_108# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_1157_298# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 a_416_86# a_452_288# a_84_108# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X17 a_27_134# a_84_108# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 a_1215_396# C a_416_86# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_1157_298# C VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X20 a_27_134# a_84_108# VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X21 VPWR A a_84_108# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
