* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 Y a_47_88# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y a_47_88# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 Y a_47_88# a_319_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_778_368# B a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_1191_368# B a_778_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 VPWR A a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 VPWR A a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_47_88# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X14 a_319_368# a_47_88# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_319_368# C a_778_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_778_368# B a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 a_319_368# C a_778_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VGND a_47_88# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 a_319_368# a_47_88# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 a_778_368# C a_319_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_778_368# C a_319_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 a_1191_368# B a_778_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_1191_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X28 a_47_88# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 VPWR D_N a_47_88# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X31 a_1191_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X32 VGND a_47_88# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 Y a_47_88# a_319_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
