* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_27_368# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_193_48# a_27_368# a_618_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VPWR a_193_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 a_892_392# A2 a_193_48# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X4 X a_193_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_193_48# A2 a_892_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 VPWR a_27_368# a_193_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 VPWR A1 a_892_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 X a_193_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 a_27_368# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 X a_193_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_618_94# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_892_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X13 a_618_94# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_618_94# a_27_368# a_193_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 VGND a_193_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_193_48# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X17 VGND A1 a_618_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 VGND a_193_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 X a_193_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VGND A2 a_618_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 VPWR a_193_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
