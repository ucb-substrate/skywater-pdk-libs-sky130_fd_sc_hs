* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
X0 VGND GATE_N a_232_98# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VGND a_27_136# a_569_79# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VGND a_647_79# a_887_270# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_27_136# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X4 VPWR a_887_270# a_1442_94# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 a_27_136# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 a_647_79# a_232_98# a_814_392# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X7 VPWR a_647_79# a_887_270# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VPWR a_27_136# a_565_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 VPWR a_887_270# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_565_392# a_343_74# a_647_79# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 Q a_887_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND a_1442_94# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 Q_N a_1442_94# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 VGND a_887_270# a_1442_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 VPWR GATE_N a_232_98# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X16 a_343_74# a_232_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_839_123# a_887_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 Q_N a_1442_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VGND a_887_270# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_343_74# a_232_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X21 a_647_79# a_343_74# a_839_123# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 Q a_887_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 a_814_392# a_887_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X24 VPWR a_1442_94# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 a_569_79# a_232_98# a_647_79# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
