* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
X0 SUM a_83_21# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 COUT a_410_58# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_1849_374# a_879_55# a_811_379# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_879_55# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_231_132# a_811_379# a_83_21# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_1660_374# a_879_55# a_1023_379# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_1023_379# B a_1849_374# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_1849_374# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_410_58# a_1023_379# a_231_132# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_1849_374# a_879_55# a_1023_379# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 a_644_104# a_811_379# a_83_21# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X11 VGND a_231_132# a_644_104# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 VGND A a_2342_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_879_55# a_811_379# a_410_58# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_1849_374# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 a_410_58# a_1023_379# a_879_55# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X16 a_83_21# a_1023_379# a_231_132# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X17 SUM a_83_21# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_811_379# B a_1660_374# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_231_132# a_811_379# a_410_58# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X20 a_83_21# a_1023_379# a_644_104# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 VPWR a_231_132# a_644_104# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X22 VPWR A a_2342_48# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X23 a_1023_379# B a_1660_374# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X24 a_1660_374# a_2342_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_1660_374# a_879_55# a_811_379# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X26 a_1660_374# a_2342_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 VPWR CI a_231_132# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X28 a_879_55# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 VGND CI a_231_132# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X30 COUT a_410_58# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 a_811_379# B a_1849_374# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
.ends
