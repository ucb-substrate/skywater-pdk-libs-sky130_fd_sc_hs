* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__clkbuf_16 A VGND VNB VPB VPWR X
X0 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X8 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_114_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_114_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 VPWR A a_114_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X28 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X30 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 VGND A a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 VPWR A a_114_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X37 VGND A a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
