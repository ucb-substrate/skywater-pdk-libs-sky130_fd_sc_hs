* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nor4bb_4 A B C_N D_N VGND VNB VPB VPWR Y
X0 a_27_368# B a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_897_349# a_864_48# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VGND a_864_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 Y a_1162_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND a_864_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_116_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_897_349# a_1162_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_27_368# a_864_48# a_897_349# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_116_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 VGND a_1162_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND D_N a_1162_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 Y a_1162_48# a_897_349# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_864_48# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X21 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 VGND a_1162_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_27_368# a_864_48# a_897_349# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 VGND C_N a_864_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_897_349# a_864_48# a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 Y a_1162_48# a_897_349# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 Y a_1162_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 VPWR D_N a_1162_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X30 a_1162_48# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X31 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 Y a_864_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 a_27_368# B a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X34 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 a_897_349# a_1162_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X36 VPWR C_N a_864_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X37 Y a_864_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
