* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nor3_4 A B C VGND VNB VPB VPWR Y
X0 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_295_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_27_368# B a_295_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 Y C a_295_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_295_368# C Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 Y C a_295_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_27_368# B a_295_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_295_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_295_368# C Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
