* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__fa_4 A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_418_74# B a_535_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 a_1141_347# B a_1235_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 VGND CIN a_734_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_734_74# a_418_74# a_1024_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR CIN a_737_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 a_737_347# a_418_74# a_1024_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 VGND A a_734_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR a_1024_74# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VPWR a_418_74# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 COUT a_418_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_737_347# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 a_1024_74# CIN a_1160_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1024_74# CIN a_1141_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X14 VPWR A a_737_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 a_1235_347# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X16 VPWR a_1024_74# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_27_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X18 COUT a_418_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 a_27_392# CIN a_418_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X20 VGND a_1024_74# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 COUT a_418_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 VGND a_418_74# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 SUM a_1024_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 a_1238_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 SUM a_1024_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 SUM a_1024_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_418_74# B a_532_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_1160_74# B a_1238_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_535_347# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X30 VPWR a_418_74# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 a_27_74# CIN a_418_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 a_532_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 VGND a_1024_74# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 VGND a_418_74# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 VPWR B a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X36 SUM a_1024_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X37 COUT a_418_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X38 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 a_734_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
