* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nand3b_1 A_N B C VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_27_116# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 a_27_116# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X4 a_269_78# B a_347_78# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND C a_269_78# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_347_78# a_27_116# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR a_27_116# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
