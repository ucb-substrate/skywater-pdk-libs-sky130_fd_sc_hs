* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_27_74# a_270_48# a_201_392# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR A2_N a_270_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 VPWR B1 a_117_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 a_500_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_270_48# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 X a_201_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 a_270_48# A2_N a_500_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_201_392# a_270_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 X a_201_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_117_392# B2 a_201_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 a_27_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND a_201_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VPWR a_201_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
