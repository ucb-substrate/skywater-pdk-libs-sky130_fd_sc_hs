* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__bufbuf_8 A VGND VNB VPB VPWR X
X0 a_27_112# A VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X1 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_334_368# a_221_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 VGND a_221_368# a_334_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_334_368# a_221_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 VPWR a_221_368# a_334_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 a_27_112# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X20 VGND a_27_112# a_221_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_334_368# a_221_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VPWR a_27_112# a_221_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 a_334_368# a_221_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
