* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__ha_2 A B VGND VNB VPB VPWR COUT SUM
X0 a_391_388# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 a_278_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_391_388# a_27_74# a_278_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VGND a_27_74# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR A a_307_388# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 VPWR a_391_388# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VPWR a_27_74# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 COUT a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 COUT a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 VPWR B a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 SUM a_391_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_307_388# B a_391_388# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X13 SUM a_391_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VGND A a_278_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VGND a_391_388# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_27_74# B a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
