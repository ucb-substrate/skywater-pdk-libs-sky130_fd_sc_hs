* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__fah_4 A B CI VGND VNB VPB VPWR COUT SUM
X0 a_1183_102# a_1378_125# VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 a_536_114# a_586_257# a_427_362# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 a_1378_125# CI VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 a_427_362# B a_536_114# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 SUM a_1278_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_586_257# a_528_362# a_1265_379# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 COUT a_1265_379# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 SUM a_1278_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VGND A a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 COUT a_1265_379# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VGND a_1265_379# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VGND a_1265_379# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_1378_125# CI VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 VPWR a_27_74# a_427_362# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_200_74# B a_528_362# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_1183_102# a_528_362# a_1278_102# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X17 a_427_362# B a_528_362# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X18 a_1278_102# a_536_114# a_1378_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_1183_102# a_1378_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_1278_102# a_536_114# a_1183_102# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X21 VGND a_27_74# a_427_362# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 VPWR a_1278_102# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 VGND B a_586_257# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 COUT a_1265_379# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_200_74# B a_536_114# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X26 VPWR B a_586_257# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 VPWR a_1265_379# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X28 a_1378_125# a_528_362# a_1265_379# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X29 SUM a_1278_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X30 a_528_362# a_586_257# a_200_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X31 a_1378_125# a_528_362# a_1278_102# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X32 VPWR a_1265_379# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X33 VPWR a_1278_102# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X34 a_1265_379# a_536_114# a_586_257# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X35 VGND a_1278_102# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 COUT a_1265_379# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X37 a_536_114# a_586_257# a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X38 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X39 VGND a_1278_102# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X40 VPWR A a_200_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X41 a_1265_379# a_536_114# a_1378_125# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X42 a_528_362# a_586_257# a_427_362# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X43 SUM a_1278_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
