* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 a_357_378# a_27_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X1 VPWR D_N a_216_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 a_357_378# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X3 VGND D_N a_216_424# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X4 a_626_378# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 a_27_424# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X6 VGND B a_357_378# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X7 a_530_378# B a_626_378# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 a_446_378# a_27_424# a_530_378# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 VPWR a_357_378# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_27_424# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X11 VGND a_216_424# a_357_378# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X12 a_357_378# a_216_424# a_446_378# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X13 VGND a_357_378# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
