* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_339_368# A4 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_788_368# A3 a_339_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_339_368# A4 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_339_368# A3 a_788_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_1191_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_1191_368# A2 a_788_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_1191_368# A2 a_788_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VPWR A1 a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_1191_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 VGND A4 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 Y A4 a_339_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_339_368# A3 a_788_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 Y A4 a_339_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 VPWR A1 a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 a_788_368# A3 a_339_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 a_27_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VGND A4 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_788_368# A2 a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X30 a_27_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 a_788_368# A2 a_1191_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X32 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
