* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__ebufn_2 A TE_B VGND VNB VPB VPWR Z
X0 VPWR TE_B a_33_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_283_48# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 VGND A a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_33_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 VPWR A a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 a_27_74# a_283_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_283_48# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 Z a_84_48# a_33_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 VGND a_283_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_33_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
