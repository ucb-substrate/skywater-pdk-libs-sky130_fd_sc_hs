* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y a_27_398# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_27_398# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 VPWR B_N a_226_398# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X3 a_435_74# a_226_398# a_513_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR a_226_398# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_627_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND B_N a_226_398# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X7 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 a_513_74# C a_627_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 Y a_27_398# a_435_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_27_398# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
.ends
