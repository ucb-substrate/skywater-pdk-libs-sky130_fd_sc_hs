* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
X0 a_1229_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 Y a_232_114# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 Y a_27_114# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 Y a_27_114# a_374_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_374_74# a_27_114# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR a_27_114# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 a_1229_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_828_74# a_232_114# a_374_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_27_114# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_374_74# a_27_114# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR a_232_114# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 VGND B_N a_232_114# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 Y a_27_114# a_374_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_1229_74# C a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 a_374_74# a_232_114# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_27_114# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X20 a_232_114# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X21 VPWR a_232_114# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 a_1229_74# C a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 a_828_74# a_232_114# a_374_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 a_828_74# C a_1229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 Y a_27_114# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X28 Y a_232_114# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X30 a_828_74# C a_1229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 VPWR A_N a_27_114# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X32 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X33 VPWR a_27_114# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X34 VGND D a_1229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 VGND D a_1229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 a_374_74# a_232_114# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 VPWR B_N a_232_114# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
.ends
