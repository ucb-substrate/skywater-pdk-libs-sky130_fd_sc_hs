* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_97_296# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_97_296# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_371_74# A2 a_449_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 X a_97_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 VPWR A3 a_362_368# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 VPWR A1 a_362_368# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 a_362_368# B1 a_97_296# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 VGND a_97_296# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND A3 a_371_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_362_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 a_449_74# A1 a_97_296# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 X a_97_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
