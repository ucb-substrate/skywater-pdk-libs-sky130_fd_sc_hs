* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
X0 VGND a_465_249# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_217_368# B a_318_389# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 VPWR A a_217_368# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 VGND A a_936_75# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_315_75# CIN a_69_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_318_389# CIN a_69_260# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 a_237_75# B a_315_75# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_69_260# a_465_249# a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VGND B a_1100_75# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 SUM a_69_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_465_249# CIN a_1100_75# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 a_509_347# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X12 VGND A a_237_75# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 VPWR A a_509_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X14 a_509_347# CIN VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 a_1107_347# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X16 VPWR a_465_249# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 VPWR B a_1107_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X18 a_1100_75# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_69_260# a_465_249# a_509_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X20 a_501_75# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 a_936_75# B a_465_249# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 a_501_75# CIN VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 VPWR A a_916_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X24 a_916_347# B a_465_249# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X25 VGND A a_501_75# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X26 a_465_249# CIN a_1107_347# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X27 SUM a_69_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
