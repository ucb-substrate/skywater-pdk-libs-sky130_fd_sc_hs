* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfxbp_1 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VPWR a_1529_74# a_1723_48# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 VPWR a_2216_94# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_1021_100# a_612_74# a_1180_496# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X3 a_233_464# D a_296_74# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X4 VPWR CLK a_612_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 VGND CLK a_612_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND a_1021_100# a_1243_398# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X7 VGND a_1723_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_218_74# D a_296_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 a_31_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X10 VGND a_31_74# a_218_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 a_2216_94# a_1723_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_434_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 a_1681_74# a_1723_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 a_1180_496# a_1243_398# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X15 a_31_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 VPWR a_1723_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 VPWR SCE a_233_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X18 a_296_74# a_828_74# a_1021_100# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X19 a_1529_74# a_828_74# a_1691_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X20 a_1243_398# a_828_74# a_1529_74# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X21 a_296_74# a_31_74# a_407_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X22 VPWR a_1021_100# a_1243_398# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X23 a_1691_508# a_1723_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X24 a_296_74# SCE a_434_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_1157_100# a_1243_398# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 VPWR a_612_74# a_828_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 a_2216_94# a_1723_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X28 a_296_74# a_612_74# a_1021_100# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 VGND a_1529_74# a_1723_48# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X30 a_1021_100# a_828_74# a_1157_100# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 a_407_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X32 VGND a_2216_94# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 VGND a_612_74# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 a_1243_398# a_612_74# a_1529_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X35 a_1529_74# a_612_74# a_1681_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
