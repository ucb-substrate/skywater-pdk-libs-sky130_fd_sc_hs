* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nor4_4 A B C D VGND VNB VPB VPWR Y
X0 Y D a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VPWR A a_879_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_496_368# C a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 VGND D Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_879_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 a_496_368# C a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 a_496_368# B a_879_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 a_879_368# B a_496_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 Y D a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_496_368# B a_879_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_27_368# C a_496_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 VPWR A a_879_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 a_27_368# C a_496_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_27_368# D Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 a_879_368# B a_496_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_879_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 Y D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_27_368# D Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
