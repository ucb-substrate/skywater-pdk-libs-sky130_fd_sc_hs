* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 X a_154_135# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VGND a_154_135# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_1102_392# C1 a_154_135# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 a_154_135# A1 a_71_135# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_1346_123# B1 a_154_135# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_1102_392# B2 a_157_376# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 VGND A2 a_71_135# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_157_376# B1 a_1102_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 X a_154_135# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 VGND B2 a_1346_123# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_157_376# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 X a_154_135# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_154_135# B1 a_1346_123# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 VGND C1 a_154_135# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_71_135# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_157_376# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X16 a_1346_123# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 a_154_135# C1 a_1102_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X18 a_1102_392# B1 a_157_376# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X19 a_154_135# C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_157_376# B2 a_1102_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X21 VPWR a_154_135# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 VPWR A2 a_157_376# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X23 VPWR a_154_135# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 X a_154_135# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VPWR A1 a_157_376# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X26 a_71_135# A1 a_154_135# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X27 VGND a_154_135# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
