* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__xor2_4 A B VGND VNB VPB VPWR X
X0 a_36_392# B a_160_98# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 a_514_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_877_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 X a_160_98# a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 a_514_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_877_74# B X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_36_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 X a_160_98# a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 a_514_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 VGND A a_877_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VGND A a_877_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 X B a_877_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 X B a_877_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_877_74# B X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR A a_36_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 VPWR A a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 a_160_98# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_160_98# B a_36_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X18 a_514_368# a_160_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 VPWR B a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 VGND A a_160_98# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VGND B a_160_98# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_514_368# a_160_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 VPWR A a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 VPWR B a_514_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 a_877_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_514_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 a_160_98# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 X a_160_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 VGND a_160_98# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
