* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=1
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=1
X2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=1
X3 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=1
.ends
