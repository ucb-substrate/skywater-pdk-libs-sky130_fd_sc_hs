* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_116_387# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 a_116_387# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 VGND a_216_387# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_27_125# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VPWR a_216_387# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_116_387# A2 a_216_387# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 VPWR B1 a_216_387# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 X a_216_387# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 X a_216_387# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND A1 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 VGND a_216_387# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VPWR a_216_387# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_216_387# B1 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_27_125# B1 a_216_387# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_27_125# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 X a_216_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 X a_216_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_216_387# A2 a_116_387# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X18 VGND A2 a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_216_387# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
.ends
