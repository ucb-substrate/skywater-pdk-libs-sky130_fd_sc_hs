* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_509_392# C1 a_148_260# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 VGND A2 a_417_79# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_310_392# B2 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 a_417_79# A1 a_148_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 X a_148_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_148_260# B1 a_597_79# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_310_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 a_509_392# B1 a_310_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 VGND C1 a_148_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 X a_148_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_597_79# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VPWR A2 a_310_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
