* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux2i_4 A0 A1 S VGND VNB VPB VPWR Y
X0 Y A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_114_85# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND a_1030_268# a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_1030_268# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 a_475_85# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_114_85# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_116_368# a_1030_268# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 Y A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 a_475_85# a_1030_268# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 Y A0 a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_478_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 VPWR S a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_475_85# A0 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1030_268# S VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X14 Y A1 a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 Y A0 a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_478_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_116_368# a_1030_268# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 a_116_368# A1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 Y A1 a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 Y A0 a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_116_368# A1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 a_114_85# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_475_85# a_1030_268# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 VPWR S a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 VGND S a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VGND S a_1030_268# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VGND a_1030_268# a_475_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_478_368# S VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 VPWR S a_1030_268# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X30 VGND S a_114_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 Y A0 a_478_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X32 a_478_368# A0 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X33 VPWR a_1030_268# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X34 a_114_85# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
