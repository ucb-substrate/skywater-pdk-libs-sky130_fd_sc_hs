* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VPWR A1 a_1330_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_1330_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 a_861_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 a_861_368# A2 a_1330_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 Y A3 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_1330_368# A2 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_27_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_27_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 a_861_368# A2 a_1330_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_1330_368# A2 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X28 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X32 a_861_368# A3 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X33 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X34 Y A3 a_861_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X35 a_27_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 VPWR A1 a_1330_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X37 a_1330_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X38 VGND A3 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
