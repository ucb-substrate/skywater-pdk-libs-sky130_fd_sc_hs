* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VPWR a_133_387# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_518_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND B2 a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR B1 a_796_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 Y B2 a_796_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_134_74# A2_N a_133_387# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VGND B1 a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_796_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VGND A1_N a_134_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_518_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR A1_N a_133_387# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X11 a_133_387# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X12 a_518_74# a_133_387# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_796_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 VPWR A2_N a_133_387# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 a_134_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 a_133_387# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X17 Y a_133_387# a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 Y a_133_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 a_133_387# A2_N a_134_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
