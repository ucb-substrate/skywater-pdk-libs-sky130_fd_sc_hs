* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1328_463# a_1369_71# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X1 VPWR a_1221_97# a_1369_71# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 a_413_90# a_850_74# a_1221_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 VGND a_1747_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VGND a_850_74# a_1023_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_850_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_413_90# SCE a_545_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 VPWR RESET_B a_2008_48# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X8 VGND a_2513_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_225_90# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 VPWR RESET_B a_413_90# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X11 a_1747_74# a_1023_74# a_1969_489# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X12 VGND RESET_B a_2124_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 a_1969_489# a_2008_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 a_1399_97# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 a_1966_74# a_2008_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 a_413_90# a_27_74# a_512_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X17 a_1321_97# a_1369_71# a_1399_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X19 a_312_90# D a_413_90# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 a_2513_424# a_1747_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X21 VPWR RESET_B a_1221_97# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X22 a_1747_74# a_850_74# a_1966_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 a_1369_71# a_850_74# a_1747_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X24 a_512_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X25 a_850_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 a_413_90# a_1023_74# a_1221_97# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X27 a_2008_48# a_1747_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X28 VPWR a_1747_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 VPWR SCE a_338_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X30 a_1221_97# a_850_74# a_1328_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X31 a_2513_424# a_1747_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X32 a_2124_74# a_1747_74# a_2008_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 a_1369_71# a_1023_74# a_1747_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X34 VPWR a_850_74# a_1023_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X35 a_545_97# SCD a_225_90# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 a_1221_97# a_1023_74# a_1321_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 VGND a_1221_97# a_1369_71# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X38 a_225_90# a_27_74# a_312_90# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 a_338_464# D a_413_90# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X40 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X41 VPWR a_2513_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
