* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VGND A3 a_351_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_330_392# B1 a_660_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 VPWR A1 a_330_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 a_351_74# A2 a_423_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_660_392# C1 a_21_270# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 a_21_270# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND C1 a_21_270# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_330_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 X a_21_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR A3 a_330_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 VGND a_21_270# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_423_74# A1 a_21_270# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR a_21_270# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 X a_21_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
