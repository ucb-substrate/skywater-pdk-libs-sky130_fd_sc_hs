* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
X0 VPWR A_N a_27_158# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X1 VPWR a_27_158# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VPWR D Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 Y a_27_158# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 a_225_74# B a_656_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 Y a_27_158# a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_656_74# B a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_656_74# C a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_1025_158# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y D VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_656_74# B a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_656_74# C a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1025_158# C a_656_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_1025_158# C a_656_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VGND D a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_27_158# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X17 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 Y a_27_158# a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VGND D a_1025_158# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 a_1025_158# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 a_225_74# a_27_158# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_27_158# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_225_74# a_27_158# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_225_74# B a_656_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
