* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__xor3_4 A B C VGND VNB VPB VPWR X
X0 a_323_392# a_397_320# a_27_118# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X1 a_1218_388# C a_416_118# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_416_118# a_1155_284# a_1218_388# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X3 a_74_294# B a_323_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X4 a_74_294# B a_416_118# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_397_320# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_323_392# a_1155_284# a_1218_388# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 X a_1218_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 a_1218_388# C a_323_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X9 VPWR a_1218_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 X a_1218_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_1155_284# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 a_27_118# a_74_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X13 a_397_320# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_1155_284# C VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X15 X a_1218_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_27_118# a_74_294# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 a_416_118# a_397_320# a_74_294# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X18 a_323_392# a_397_320# a_74_294# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 VGND A a_74_294# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 X a_1218_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VPWR A a_74_294# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X22 a_27_118# B a_323_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 VPWR a_1218_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 VGND a_1218_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_416_118# a_397_320# a_27_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 VGND a_1218_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_27_118# B a_416_118# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
.ends
