* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_1457_508# a_1470_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X1 a_1027_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 a_709_463# a_760_395# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X3 VGND a_1902_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_27_74# a_398_74# a_604_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X5 a_1215_74# a_398_74# a_1298_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_1500_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_1902_74# a_1298_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X8 a_760_395# a_604_74# a_1027_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 a_1902_74# a_1298_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 a_27_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 a_1298_392# a_398_74# a_1457_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X12 VPWR a_224_350# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_604_74# a_224_350# a_709_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 VPWR SET_B a_1298_392# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X15 VPWR a_604_74# a_1197_341# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X16 a_604_74# a_398_74# a_740_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_1422_74# a_1470_48# a_1500_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 VGND a_224_350# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VPWR a_1902_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 a_1298_392# a_224_350# a_1422_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 VGND a_604_74# a_1215_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 a_1197_341# a_224_350# a_1298_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X23 a_224_350# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_27_74# a_224_350# a_604_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 VGND a_1298_392# a_1470_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 a_224_350# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 VPWR a_604_74# a_760_395# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X28 VPWR a_1298_392# a_1470_48# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X29 a_740_74# a_760_395# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X30 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 a_760_395# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends
