* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VGND A2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND A2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 Y C1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_27_84# B1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_483_74# B1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_483_74# B2 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_483_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR B1 a_508_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 a_483_74# B1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 Y A2 a_1288_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 Y B2 a_508_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 Y A2 a_1288_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_27_84# B2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 a_508_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 VPWR A1 a_1288_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_1288_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 a_27_84# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 Y B2 a_508_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 a_483_74# B2 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_483_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_483_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VPWR A1 a_1288_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 a_1288_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 a_27_84# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_508_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 VPWR B1 a_508_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X30 a_1288_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 a_508_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X32 a_508_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X33 Y C1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 VGND A1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 VGND A1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 a_1288_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X37 a_27_84# B2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 a_27_84# B1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 a_483_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
