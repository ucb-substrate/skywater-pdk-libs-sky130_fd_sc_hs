* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 X a_137_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR A2 a_1013_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 a_137_260# D1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND A2 a_1210_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_137_260# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 X a_137_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 a_549_392# C1 a_814_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 X a_137_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 a_1013_392# B1 a_814_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 a_1013_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 a_1013_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 X a_137_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND a_137_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_137_260# A1 a_1210_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 VGND C1 a_137_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_549_392# D1 a_137_260# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X16 a_1210_74# A1 a_137_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 VPWR a_137_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 a_137_260# D1 a_549_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X19 VGND a_137_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VGND D1 a_137_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 VPWR a_137_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 a_814_392# C1 a_549_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X23 a_1210_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 VGND B1 a_137_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X25 a_814_392# B1 a_1013_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X26 a_137_260# C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X27 VPWR A1 a_1013_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
