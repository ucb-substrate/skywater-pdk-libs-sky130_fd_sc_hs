* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__bufinv_8 A VGND VNB VPB VPWR Y
X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VPWR a_27_368# a_183_48# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_183_48# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 Y a_183_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR a_183_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 Y a_183_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR a_27_368# a_183_48# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 VPWR a_183_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR a_183_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 VPWR a_183_48# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 Y a_183_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND a_27_368# a_183_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VGND a_27_368# a_183_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 Y a_183_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 a_183_48# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 Y a_183_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 VGND a_183_48# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
