* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__maj3_1 A B C VGND VNB VPB VPWR X
X0 a_223_120# B a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_226_384# B a_84_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 a_406_384# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 X a_84_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VGND A a_223_120# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_403_136# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VPWR A a_226_384# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 a_595_136# C a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_84_74# B a_406_384# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 a_598_384# C a_84_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 VGND A a_595_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 X a_84_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_84_74# B a_403_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 VPWR A a_598_384# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
