* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__fah_2 A B CI VGND VNB VPB VPWR COUT SUM
X0 a_1689_424# a_849_424# a_1895_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_849_424# a_481_379# a_413_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_1689_424# a_514_424# a_1895_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X3 VPWR a_1451_424# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 a_413_392# a_481_379# a_514_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X5 a_1895_424# a_849_424# a_2052_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 VPWR a_1895_424# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VGND CI a_1689_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_1451_424# a_849_424# a_1689_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X9 a_114_368# B a_849_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_114_368# a_481_379# a_849_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X11 a_481_379# a_514_424# a_1451_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X12 SUM a_1895_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 VPWR a_81_260# a_114_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 VGND A a_413_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 VGND B a_481_379# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 SUM a_1895_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_81_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 VGND a_1895_424# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_1895_424# a_514_424# a_2052_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_481_379# a_849_424# a_1451_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 a_2052_424# a_1689_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X22 VPWR A a_413_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X23 a_413_392# B a_514_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 VPWR CI a_1689_424# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X25 COUT a_1451_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 COUT a_1451_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_514_424# B a_114_368# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X28 VGND a_81_260# a_114_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_849_424# B a_413_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X30 VPWR B a_481_379# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 VGND a_1451_424# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 a_1451_424# a_514_424# a_1689_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X33 a_2052_424# a_1689_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X34 a_81_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X35 a_514_424# a_481_379# a_114_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
