* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__einvn_8 A TE_B VGND VNB VPB VPWR Z
X0 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VPWR TE_B a_126_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VGND TE_B a_126_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X28 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X30 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X33 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
