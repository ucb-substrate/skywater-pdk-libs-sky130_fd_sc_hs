* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlymetal6s4s_1 A VGND VNB VPB VPWR X
X0 VGND a_28_138# a_209_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_316_138# a_209_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 VGND a_604_138# a_785_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_28_138# a_209_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 VPWR a_316_138# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_604_138# X VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X6 VPWR a_604_138# a_785_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 a_28_138# A VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X8 VGND a_316_138# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_28_138# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 a_316_138# a_209_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 a_604_138# X VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
