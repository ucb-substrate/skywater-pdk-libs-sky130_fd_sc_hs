* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
