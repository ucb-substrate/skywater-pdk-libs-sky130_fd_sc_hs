* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_131_74# B1 a_209_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_209_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_209_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND A3 a_209_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VPWR B1 a_31_387# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 VPWR a_31_387# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 a_31_387# A3 a_320_387# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 a_536_387# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 VGND a_31_387# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_320_387# A2 a_536_387# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 a_31_387# C1 a_131_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 a_31_387# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
