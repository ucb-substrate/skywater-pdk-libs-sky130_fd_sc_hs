* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_131_383# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X1 a_490_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VPWR a_131_383# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 a_397_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y B2 a_490_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 Y a_131_383# a_397_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND B1 a_397_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR A1_N a_131_383# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X8 VGND A1_N a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_114_74# A2_N a_131_383# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
