* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VGND A3 a_264_120# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_89_270# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_359_123# A1 a_89_270# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VPWR A1 a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X4 a_264_120# A2 a_359_123# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 X a_89_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 VPWR A3 a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 X a_89_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_546_392# C1 a_89_270# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 VGND C1 a_89_270# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_258_392# B1 a_546_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 a_258_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
