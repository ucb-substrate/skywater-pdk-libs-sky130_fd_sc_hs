* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X
X0 a_355_368# a_194_125# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 X a_194_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VPWR A a_158_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 VGND A a_194_125# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X4 a_194_125# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X5 a_355_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 a_455_87# B X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR B a_355_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VGND A a_455_87# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_158_392# B a_194_125# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
