* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_452_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_1814_48# a_1587_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 a_1587_74# a_630_74# a_1766_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_301_74# SCE a_452_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_301_74# a_630_74# a_1026_100# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 Q a_1814_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_36_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 VPWR a_630_74# a_828_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 VPWR a_1026_100# a_1257_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X9 a_301_74# a_36_74# a_412_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X10 VPWR a_1814_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_1814_48# a_1587_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_36_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X13 a_1257_74# a_630_74# a_1587_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X14 VGND a_1814_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 a_1026_100# a_630_74# a_1214_506# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X16 Q a_1814_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 VGND a_1026_100# a_1257_74# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X18 a_1026_100# a_828_74# a_1162_100# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 a_1162_100# a_1257_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 a_1257_74# a_828_74# a_1587_74# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X21 a_412_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X22 VPWR SCE a_238_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X23 a_1214_506# a_1257_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X24 VPWR CLK a_630_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 VGND a_1814_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VPWR a_1587_74# a_1814_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X27 a_238_464# D a_301_74# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X28 a_1587_74# a_828_74# a_1764_476# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X29 VGND CLK a_630_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 Q a_1814_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 a_301_74# a_828_74# a_1026_100# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X32 a_1764_476# a_1814_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X33 VPWR a_1814_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X34 a_223_74# D a_301_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 Q a_1814_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 VGND a_36_74# a_223_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 VGND a_630_74# a_828_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 a_1766_74# a_1814_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
