* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 VPWR a_1338_125# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_846_74# S0 a_979_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_1338_125# a_1396_99# a_342_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_1396_99# S1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_255_341# S0 a_342_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 a_264_74# a_27_74# a_342_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_846_74# S1 a_1338_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 VGND A0 a_264_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_342_74# S0 a_450_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_979_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_27_74# S0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 a_537_341# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X12 a_768_74# a_27_74# a_846_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_846_74# a_27_74# a_1065_387# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X14 a_342_74# S1 a_1338_125# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 VGND a_1338_125# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND A2 a_768_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 a_1065_387# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X18 a_342_74# a_27_74# a_537_341# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X19 a_450_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_763_341# S0 a_846_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X21 VPWR A0 a_255_341# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X22 a_1338_125# a_1396_99# a_846_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X23 a_1396_99# S1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X24 VPWR A2 a_763_341# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X25 a_27_74# S0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
