* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__xnor2_2 A B VGND VNB VPB VPWR Y
X0 VGND A a_340_107# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 Y B a_638_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_151_74# B a_133_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_340_107# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y a_133_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_638_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 Y a_133_368# a_340_107# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR A a_133_368# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 a_340_107# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND B a_340_107# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR A a_638_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_638_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 VPWR a_133_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_133_368# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X14 VGND A a_151_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 a_340_107# a_133_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
