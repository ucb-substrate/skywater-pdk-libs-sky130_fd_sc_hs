* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_510_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 Y A2 a_697_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 VGND A2 a_510_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_299_74# B1 a_510_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND A1 a_510_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR A1 a_697_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 a_510_74# B1 a_299_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_510_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_697_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_299_74# C1 a_40_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_697_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_40_74# D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 a_40_74# C1 a_299_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 Y D1 a_40_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
