* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__ebufn_8 A TE_B VGND VNB VPB VPWR Z
X0 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_833_48# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 a_27_74# a_833_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 VGND A a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 Z a_84_48# a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 Z a_84_48# a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 VPWR A a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 Z a_84_48# a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 a_84_48# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 Z a_84_48# a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 a_27_74# a_833_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_28_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 VPWR TE_B a_28_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 VGND a_833_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_27_74# a_833_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_27_74# a_833_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_28_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 VGND a_833_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_28_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X28 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_84_48# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 a_28_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 Z a_84_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 VGND a_833_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 a_833_48# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 a_27_74# a_84_48# Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 a_28_368# a_84_48# Z VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X37 VGND a_833_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
