* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_95_306# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VGND A2 a_1064_123# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_1064_123# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_555_392# B2 a_95_306# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X4 a_95_306# B2 a_555_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 a_95_306# B1 a_645_120# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VPWR a_95_306# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 a_1064_123# A1 a_95_306# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_95_306# A1 a_1064_123# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 VPWR A1 a_555_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 a_555_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 VGND a_95_306# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR a_95_306# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 VGND B2 a_645_120# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_95_306# B1 a_555_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 VGND a_95_306# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_555_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X17 X a_95_306# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_645_120# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_555_392# B1 a_95_306# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X20 a_645_120# B1 a_95_306# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 X a_95_306# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 X a_95_306# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 VPWR A2 a_555_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
