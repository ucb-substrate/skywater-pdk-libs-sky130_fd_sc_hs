* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A2 a_71_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_71_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 Y A1 a_339_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_339_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_159_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_71_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 Y B1 a_71_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VGND B2 a_159_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
