* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VPWR a_194_136# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_34_392# a_272_110# a_194_136# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 VGND a_194_136# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_194_136# a_272_110# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_122_136# A1 a_194_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_34_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 a_272_110# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 VPWR A1 a_34_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 VGND A2 a_122_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_272_110# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
.ends
