* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a222o_2 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
X0 a_639_368# B1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 a_27_82# C1 a_114_82# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_775_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND a_27_82# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_27_82# B1 a_775_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 X a_27_82# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 X a_27_82# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND A2 a_557_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_27_82# C1 a_116_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 VPWR A1 a_639_368# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 a_639_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 a_116_392# B2 a_639_368# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X12 VPWR a_27_82# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_557_74# A1 a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_116_392# C2 a_27_82# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 a_114_82# C2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
