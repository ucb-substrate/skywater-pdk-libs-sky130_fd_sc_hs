* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_491_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR a_81_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 a_81_48# B2 a_388_368# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 a_388_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X4 X a_81_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VPWR A1 a_388_368# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X6 VGND a_81_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_81_48# B1 a_491_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_304_74# A1 a_81_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 X a_81_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X10 VGND A2 a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_388_368# B1 a_81_48# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
