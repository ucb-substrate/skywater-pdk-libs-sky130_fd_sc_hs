* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_83_244# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 a_651_78# B1 a_564_78# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 X a_83_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 VGND a_83_244# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR A1 a_1338_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 VGND A3 a_564_78# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_564_78# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_564_78# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_83_244# C1 a_651_78# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 VGND A1 a_564_78# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 VPWR B1 a_83_244# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 VGND a_83_244# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR C1 a_83_244# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X13 a_83_244# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X14 a_83_244# A3 a_1034_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 a_651_78# C1 a_83_244# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 X a_83_244# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_1338_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X18 VGND A2 a_564_78# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_83_244# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X20 X a_83_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 a_564_78# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 a_1034_392# A3 a_83_244# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X23 VPWR a_83_244# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 a_1034_392# A2 a_1338_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X25 X a_83_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_1338_392# A2 a_1034_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X27 a_564_78# B1 a_651_78# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
