* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__ha_4 A B VGND VNB VPB VPWR COUT SUM
X0 SUM a_294_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR B a_435_99# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 VGND B a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_435_99# A VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X4 COUT a_435_99# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_707_119# B a_435_99# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 SUM a_294_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 a_294_392# a_435_99# a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VGND a_435_99# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND a_294_392# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR A a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 a_435_99# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X12 VGND a_294_392# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_294_392# B a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X14 SUM a_294_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 VGND a_435_99# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_294_392# a_435_99# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X17 a_435_99# B a_707_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 COUT a_435_99# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 SUM a_294_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 COUT a_435_99# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_27_125# a_435_99# a_294_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 VGND A a_707_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 a_27_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 VPWR a_435_99# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 a_27_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X26 a_707_119# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X27 COUT a_435_99# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 VPWR a_294_392# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 a_27_125# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X30 VPWR a_294_392# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 a_27_392# B a_294_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X32 VPWR A a_435_99# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X33 VGND A a_27_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X34 VPWR a_435_99# a_294_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X35 VPWR a_435_99# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
