* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__or3_4 A B C VGND VNB VPB VPWR X
X0 X a_302_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_206_388# C a_302_388# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X2 a_116_388# B a_206_388# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 VGND B a_302_388# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_302_388# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 X a_302_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 X a_302_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VPWR A a_116_388# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 a_302_388# C a_206_388# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 a_206_388# B a_116_388# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 a_302_388# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 X a_302_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND a_302_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VPWR a_302_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_116_388# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 VPWR a_302_388# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 VGND a_302_388# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
