* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_27_79# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_2158_74# a_1790_74# a_2006_373# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 VGND a_2604_392# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_1323_118# a_1370_289# a_1401_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_307_464# D a_388_79# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X5 a_223_79# a_27_79# a_310_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_388_79# a_27_79# a_538_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X7 a_388_79# SCE a_547_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X8 VPWR a_2604_392# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 a_223_79# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 VPWR a_1223_118# a_1370_289# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 a_388_79# a_852_74# a_1223_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 VGND RESET_B a_2158_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 VGND a_1790_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 Q a_2604_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VGND a_1790_74# a_2604_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 a_538_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X17 Q_N a_1790_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 a_1401_118# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 a_2000_74# a_2006_373# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 VPWR SCE a_307_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X21 a_2006_373# a_1790_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X22 a_388_79# a_1025_74# a_1223_118# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X23 a_1223_118# a_1025_74# a_1323_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 a_1223_118# a_852_74# a_1325_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X25 a_1790_74# a_852_74# a_2000_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 a_852_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 VGND a_1223_118# a_1370_289# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X28 a_310_79# D a_388_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 VPWR a_1790_74# a_2604_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X30 Q a_2604_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 VPWR a_852_74# a_1025_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X32 a_1325_457# a_1370_289# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X33 a_1955_471# a_2006_373# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X34 a_27_79# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X35 a_1370_289# a_852_74# a_1790_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X36 VPWR a_1790_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X37 a_547_79# SCD a_223_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 VPWR RESET_B a_1223_118# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X39 VGND a_852_74# a_1025_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X40 a_1790_74# a_1025_74# a_1955_471# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X41 a_852_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X42 VPWR RESET_B a_2006_373# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X43 Q_N a_1790_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X44 a_1370_289# a_1025_74# a_1790_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X45 VPWR RESET_B a_388_79# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
.ends
