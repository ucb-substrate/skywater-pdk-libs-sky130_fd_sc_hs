* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VGND A1 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_132_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_132_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_314_368# A4 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_314_368# A3 a_607_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 a_607_368# A2 a_807_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X8 Y B1 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_132_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_807_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 VGND A2 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 Y A4 a_314_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_607_368# A3 a_314_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_807_368# A2 a_607_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 a_132_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND A4 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VGND A3 a_132_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_132_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VPWR A1 a_807_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
