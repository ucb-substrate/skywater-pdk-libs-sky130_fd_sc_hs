* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
X0 VGND CLK_N a_300_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VPWR a_300_74# a_507_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VPWR D a_33_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X3 a_120_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_714_127# a_300_74# a_850_127# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 a_1550_119# a_1598_93# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 VPWR RESET_B a_1598_93# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X7 a_1598_93# a_1266_119# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X8 a_714_127# a_507_368# a_817_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X9 VPWR RESET_B a_714_127# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X10 a_1266_119# a_507_368# a_1550_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 VGND a_714_127# a_856_304# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_33_74# D a_120_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 a_1547_508# a_1598_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 a_33_74# a_507_368# a_714_127# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 a_817_508# a_856_304# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X16 VGND RESET_B a_1736_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_850_127# a_856_304# a_922_127# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 a_922_127# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 a_1934_94# a_1266_119# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X20 VPWR a_1934_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_1736_119# a_1266_119# a_1598_93# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 a_33_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X23 a_33_74# a_300_74# a_714_127# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X24 a_856_304# a_300_74# a_1266_119# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VPWR CLK_N a_300_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X26 a_856_304# a_507_368# a_1266_119# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X27 a_1934_94# a_1266_119# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X28 VGND a_1934_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 VGND a_300_74# a_507_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 VPWR a_714_127# a_856_304# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X31 a_1266_119# a_300_74# a_1547_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends
