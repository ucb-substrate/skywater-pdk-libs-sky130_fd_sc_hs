* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__bufinv_16 A VGND VNB VPB VPWR Y
X0 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X2 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VGND a_27_74# a_384_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X19 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X23 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X24 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 VPWR a_27_74# a_384_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X29 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X30 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 Y a_384_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X33 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X34 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X35 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X37 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X38 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X39 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X40 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X41 VPWR a_384_74# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X42 a_384_74# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X43 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X44 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X45 a_384_74# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X46 Y a_384_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X47 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X48 VGND a_384_74# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X49 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
