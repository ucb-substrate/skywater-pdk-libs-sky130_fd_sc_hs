* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 VPWR a_998_81# a_1610_341# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 a_1721_374# a_1958_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X2 a_2395_94# a_1764_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_1128_457# a_1198_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X4 a_599_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND a_2395_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_1764_74# a_599_74# a_1610_341# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 a_1686_74# a_800_74# a_1764_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_238_74# D a_289_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 a_998_81# a_800_74# a_1150_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 VGND a_998_81# a_1686_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VPWR a_2395_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X12 a_1910_74# a_1958_48# a_1988_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 a_1426_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 a_1988_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 a_402_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 a_1958_48# a_1764_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X17 VPWR a_599_74# a_800_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X18 a_998_81# a_599_74# a_1128_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X19 a_289_464# SCE a_402_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 a_289_464# a_599_74# a_998_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 VPWR SCE a_205_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X22 a_2395_94# a_1764_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X23 VGND a_27_464# a_238_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 a_1150_81# a_1198_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_289_464# a_27_464# a_415_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X26 VPWR SET_B a_1764_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X27 a_205_464# D a_289_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X28 VGND a_1764_74# a_1958_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 a_1198_55# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X30 a_1721_374# a_800_74# a_1764_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X31 a_289_464# a_800_74# a_998_81# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X32 a_1764_74# a_599_74# a_1910_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 a_415_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X34 VPWR a_998_81# a_1198_55# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X35 a_1198_55# a_998_81# a_1426_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 VGND a_599_74# a_800_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 a_27_464# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 a_27_464# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X39 a_599_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
.ends
