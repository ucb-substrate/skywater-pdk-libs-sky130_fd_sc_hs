* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_83_283# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X1 VGND a_83_283# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_83_283# B1 a_587_110# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND A3 a_992_122# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VPWR A1 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X5 VGND a_83_283# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_587_110# B1 a_83_283# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_1079_122# A2 a_992_122# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_509_392# B1 a_83_283# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 a_509_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 X a_83_283# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_992_122# A2 a_1079_122# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_587_110# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 X a_83_283# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_83_283# B2 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X15 VPWR A3 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X16 a_509_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X17 a_1079_122# A1 a_83_283# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 a_992_122# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 X a_83_283# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 VPWR A2 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X21 a_509_392# B2 a_83_283# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X22 a_83_283# A1 a_1079_122# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 VGND B2 a_587_110# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 VPWR a_83_283# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 a_509_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X26 X a_83_283# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_83_283# B1 a_509_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
.ends
