* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 VGND RESET_B a_1624_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_125_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 VPWR a_1224_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 a_38_78# D a_125_78# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 VGND a_319_360# a_498_360# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_910_118# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 VPWR a_319_360# a_498_360# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VGND a_1224_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR a_706_463# a_841_401# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 a_841_401# a_319_360# a_1224_74# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X10 a_1434_74# a_1482_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 a_1224_74# a_498_360# a_1465_471# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X12 VPWR a_2026_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_706_463# a_319_360# a_796_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 VPWR RESET_B a_706_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X15 a_1482_48# a_1224_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X16 a_38_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X17 a_1465_471# a_1482_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X18 VGND a_2026_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_319_360# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_2026_424# a_1224_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X21 a_38_78# a_319_360# a_706_463# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 a_796_463# a_841_401# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X23 VGND a_706_463# a_841_401# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 a_319_360# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X25 a_1224_74# a_319_360# a_1434_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 a_2026_424# a_1224_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X27 a_706_463# a_498_360# a_832_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X28 a_841_401# a_498_360# a_1224_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X29 a_1624_74# a_1224_74# a_1482_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X30 VPWR D a_38_78# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X31 a_38_78# a_498_360# a_706_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X32 VPWR RESET_B a_1482_48# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X33 a_832_118# a_841_401# a_910_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
