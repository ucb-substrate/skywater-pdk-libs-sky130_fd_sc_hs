* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_615_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VGND a_212_102# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 Y a_212_102# a_424_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 Y B2 a_615_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR B2 a_424_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 VPWR B1 a_424_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X6 VPWR A1_N a_209_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X7 VGND B1 a_615_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 Y a_212_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_615_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_209_392# A2_N a_212_102# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X11 a_212_102# A2_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_424_368# a_212_102# Y VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X13 a_424_368# B2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X14 a_424_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 VGND A1_N a_212_102# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
