* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1517_508# a_1510_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X1 a_1462_74# a_1510_48# a_1540_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 a_1355_377# a_225_74# a_1462_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_779_380# a_596_81# a_1061_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_2113_74# a_1355_377# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X5 VGND a_1355_377# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_27_80# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_1355_377# a_398_74# a_1517_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X8 a_225_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X9 a_748_81# a_779_380# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 VPWR a_2113_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 a_1540_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 VPWR a_596_81# a_779_380# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X13 a_1510_48# a_1355_377# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 VPWR SET_B a_1355_377# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X15 a_2113_74# a_1355_377# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X16 VPWR a_1355_377# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 a_728_463# a_779_380# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X18 VGND a_2113_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VPWR a_596_81# a_1254_341# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X20 VGND a_596_81# a_1262_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 VGND a_225_74# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_1262_74# a_398_74# a_1355_377# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 a_27_80# a_398_74# a_596_81# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X24 a_27_80# a_225_74# a_596_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_1254_341# a_225_74# a_1355_377# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X26 a_596_81# a_398_74# a_748_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 a_225_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_1061_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 a_779_380# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X30 VPWR a_225_74# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X31 a_596_81# a_225_74# a_728_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X32 VGND a_1355_377# a_1510_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 a_27_80# D VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends
