* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_1047_74# a_27_74# a_1044_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_524_508# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X2 GCLK a_1044_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X3 a_334_54# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_27_74# a_84_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 VGND a_1044_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_1044_368# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X7 VPWR GATE a_283_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X8 VGND CLK a_1047_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 GCLK a_1044_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR CLK a_1044_368# VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X11 GCLK a_1044_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND a_1044_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_283_392# a_334_338# a_84_48# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X14 a_286_80# a_334_54# a_84_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 VPWR a_1044_368# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X16 VGND a_334_54# a_334_338# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VGND GATE a_286_80# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 VPWR a_334_54# a_334_338# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X19 GCLK a_1044_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X20 VPWR a_1044_368# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X21 a_334_54# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X22 a_491_124# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 a_84_48# a_334_54# a_524_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X24 a_27_74# a_84_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_84_48# a_334_338# a_491_124# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
