* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_27_392# A2 a_747_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X1 a_27_74# C1 a_287_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_747_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X3 VPWR C1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X4 VPWR a_27_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X5 a_27_392# D1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND a_27_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 X a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_747_392# A2 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X9 a_287_74# C1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_287_74# B1 a_477_198# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_477_198# B1 a_287_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR D1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X13 a_27_392# D1 VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X14 X a_27_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X15 VPWR B1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X16 X a_27_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X17 VPWR A1 a_747_392# VPB sky130_fd_pr__pfet_01v8 w=1 l=150000u
X18 a_477_198# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VGND A1 a_477_198# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VGND a_27_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VGND A2 a_477_198# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 X a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_477_198# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_27_74# D1 a_27_392# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_27_392# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X26 VPWR a_27_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12 l=150000u
X27 a_27_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
.ends
